45nm XOR Gate
.lib '/class/ece482/gpdk045_mos' TT

c1 vdd vss 368.19e-18
c2 a vss 248.239e-18
c3 b vss 191.528e-18
c4 f vss 139.07e-18
c5 net1 vss 148.388e-18
mpm0 f b a vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mpm1 net1 a vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mnm1 f b net1 vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm0 net1 a vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1

vSupply vdd 0 1.1
vGnd vss 0 0
vA a 0 pulse (0 1.1 0 100p 100p 2n 4n)
vB b 0 pulse (0 1.1 1n 100p 100p 2n 4n)

.tran 1p 16n
.option post
.END
