45nm XOR Gate
.lib '/class/ece482/gpdk045_mos' TT

c1 vdd vss 621.026e-18
c2 a vss 259.928e-18
c3 b vss 206.149e-18
c4 f vss 146.558e-18
c5 net2 vss 306.996e-18
c6 net1 vss 220.371e-18
mpm0 net2 b net1 vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mpm2 f net2 vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mpm1 net1 a vdd vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mnm2 net2 b a vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm3 f net2 vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm1 net1 a vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1

vSupply vdd 0 1.1
vGnd vss 0 0
vA a 0 pulse (0 1.1 0 100p 100p 2n 4n)
vB b 0 pulse (0 1.1 1n 100p 100p 2n 4n)

.tran 1p 16n
.option post
.END
